`ifndef FIFO_DEFINE_SV
`define FIFO_DEFINE_SV

`define DEPTH 16 //Depth of FIFO 
`define ADDR 4 //Address width 
`define WIDTH 8 //Data width 

`endif 

